acl:att
acl:av
acl:cleft
acl:efter
acl:från
acl:för
acl:hos
acl:i
acl:liksom
acl:med
acl:mot
acl:när
acl:om
acl:på
acl:relcl
acl:som
acl:såsom
acl:till
acl:utan
acl:vid
acl:än
acl:över
advcl:allt_efter_som
advcl:allt_eftersom
advcl:alltefter_som
advcl:allteftersom
advcl:antingen
advcl:att
advcl:av
advcl:av:om
advcl:därför_att
advcl:då
advcl:efter
advcl:efter_hand_som
advcl:eftersom
advcl:ehuruväl
advcl:emedan
advcl:fast
advcl:fastän
advcl:från
advcl:från_det
advcl:för
advcl:för_att
advcl:förrän
advcl:förutsatt_att
advcl:hos
advcl:i
advcl:innan
advcl:liksom
advcl:låt_vara
advcl:med
advcl:med:att
advcl:medan
advcl:när
advcl:nära
advcl:oavsett
advcl:oberoende_av
advcl:om
advcl:på
advcl:på:att
advcl:på_det
advcl:samtidigt_som
advcl:sedan
advcl:som
advcl:så_att
advcl:såsom
advcl:såvida
advcl:till
advcl:tills
advcl:trots_att
advcl:utan
advcl:vare_sig
advcl:än
advcl:även_om
advcl:över
aux:pass
compound:prt
conj:eller
conj:fast
conj:för
conj:men
conj:och
conj:plus
conj:resp
conj:respektive
conj:samt
conj:som
conj:såväl:som
conj:ty
conj:utan
csubj:pass
flat:name
nmod:angående
nmod:av
nmod:bak
nmod:bakom
nmod:beträffande
nmod:bland
nmod:efter
nmod:emellan
nmod:enligt
nmod:framför
nmod:från
nmod:från_och_med
nmod:för
nmod:för:i
nmod:före
nmod:genom
nmod:gentemot
nmod:hos
nmod:i
nmod:i_form_av
nmod:i_samband_med
nmod:inför
nmod:inklusive
nmod:inom
nmod:intill
nmod:jämte
nmod:kontra
nmod:kring
nmod:längs
nmod:med
nmod:med_hänsyn_till
nmod:mellan
nmod:mot
nmod:oavsett
nmod:om
nmod:omkring
nmod:ovanför
nmod:ovanpå
nmod:per
nmod:plus
nmod:poss
nmod:på
nmod:på:för
nmod:runt
nmod:rörande
nmod:sedan
nmod:till
nmod:till_och_med
nmod:trots
nmod:under
nmod:ur
nmod:utan
nmod:utanför
nmod:utom
nmod:utom:om
nmod:utöver
nmod:via
nmod:vid
nmod:än
nmod:än:med
nmod:å
nmod:åt
nmod:över
nsubj:pass
obl:agent
obl:allt_efter
obl:alltefter
obl:av
obl:bakom
obl:beträffande
obl:bland
obl:bortsett_från
obl:efter
obl:emellan
obl:enligt
obl:exklusive
obl:framemot
obl:framför
obl:från
obl:från_och_med
obl:frånsett
obl:för
obl:för_sedan
obl:för_sen
obl:för_skull
obl:före
obl:förutan
obl:förutom
obl:genom
obl:gentemot
obl:hos
obl:i
obl:i_enlighet_med
obl:i_form_av
obl:i_fråga_om
obl:i_närheten_av
obl:i_och_med
obl:i_riktning_mot
obl:i_samband_med
obl:ifråga_om
obl:ifrån
obl:igenom
obl:inför
obl:innanför
obl:inom
obl:inpå
obl:intill
obl:jämfört_med
obl:kring
obl:längs
obl:med
obl:med_avseende_på
obl:med_hänsyn_till
obl:mellan
obl:mot
obl:nedanför
obl:nedom
obl:när_det_gäller
obl:när_det_gällt
obl:nära
obl:närmare
obl:oavsett
obl:oberoende_av
obl:om
obl:omkring
obl:ovanför
obl:ovanpå
obl:per
obl:på
obl:på:till
obl:på_grund_av
obl:runtomkring
obl:sedan
obl:senast
obl:som
obl:tack_vare
obl:tidigast
obl:till
obl:till_och_med
obl:to
obl:trots
obl:tvärsigenom
obl:tvärtemot
obl:under
obl:ur
obl:utan
obl:utanför
obl:utifrån
obl:utom
obl:utåt
obl:utöver
obl:vad_beträffar
obl:via
obl:vid
obl:vid_sidan_av
obl:än
obl:å
obl:åt
obl:över
